`timescale 1ns/1ps
// Module inspired by fpu_apb_wrapper.v
module adc_apb_wrapper #(
    parameter ADDR_WIDTH = 12,
    parameter DATA_WIDTH = 32
)
(
    // Clock and reset signals
    // Clock signal which synchronises bus operations
    input  wire                  PCLK, 
    // Active-low reset signal, used to initialise bus peripherals.
    input  wire                  PRESETn,

    // Address and control signals
    // Peripheral select. There is one of these wires for every peripheral on the bus.
    input  wire                  PSEL,
    // Address bus that specifies peripheral memory location
    input  wire [ADDR_WIDTH-1:0] PADDR,
    // Indicates start of accessing phase. 
    input  wire                  PENABLE,
    // Indicates direction of data transfer. High is a write, low is read.
    input  wire                  PWRITE,

    // Data Signals
    // Write data bus. Carries data from master to peripheral during write transaction.
    input  wire [DATA_WIDTH-1:0] PWDATA,
    // Read data bus. Peripheral places data on bus during read transaction.
    output reg  [DATA_WIDTH-1:0] PRDATA,
    // Handshake signals
    // Slave indicates ready to complete data transfer.
    output reg                   PREADY,
    // Signal that indicates if an error occured during transaction.
    output wire                  PSLVERR,

    // ADC interface 
    input  wire [55:0]           adc_data,
    input  wire                  adc_data_valid
);

    // --------------------------------------------------------------------------
    // ADC wires - Connect from read and write to the actual ADC.
    // --------------------------------------------------------------------------
    // THE fpu_apb_wrapper gives an example of using this to write to the correct item.
    // This should be implemented.
    // Consider what actual inputs and outputs are needed.
    reg [DATA_WIDTH-1:0] pll_reg;
    reg [DATA_WIDTH-1:0] amux_reg;
    reg [DATA_WIDTH-1:0] trig_reg;
    // Statis_reg is used to reflect the FIFO status and ADC data validity
    reg [DATA_WIDTH-1:0] status_reg;

    // Signal used to trigger FIFO reset (generated by ADC triggering write operation)
    reg                  adc_trig;

    // FIFO signal
    wire                 fifo_full, fifo_empty;
    wire [55:0]          fifo_data_out;
    reg                  fifo_rd_en;   // Used to trigger FIFO read out
    reg                  fifo_rd_en_d; // Delay one clock cycle of Fifo'rd_den

    // --------------------------------------------------------------------------
    // APB addresses for various ADC functionality
    // --------------------------------------------------------------------------
    // These are address offsets (base + offset)
    // ADC Reads
    localparam STATUS_REG_ADDR     = 12'h001;
    localparam MEASUREMENT_HI_ADDR = 12'h002;
    localparam MEASUREMENT_LO_ADDR = 12'h003;
    // ADC Writes
    localparam PLL_CONTROL_ADDR    = 12'h100;
    localparam AMUX_ADDR           = 12'h101;
    localparam ADC_TRIGGER_ADDR    = 12'h102;

    // --------------------------------------------------------------------------
    // APB control signals
    // --------------------------------------------------------------------------
    wire read_enable  = PSEL & ~PWRITE;
    wire write_enable = PSEL & PWRITE & PENABLE;

    // --------------------------------------------------------------------------
    // Instantiate FIFO module
    // --------------------------------------------------------------------------
    fifo_apb_adc fifo (
        .clk          (PCLK),
        .rst_n        (PRESETn),
        .adc_wr_en    (adc_data_valid & ~fifo_full),
        .adc_data     (adc_data),
        .fifo_full    (fifo_full),
        .apb_rd_en    (fifo_rd_en),
        .apb_rd_data  (fifo_data_out),
        .fifo_empty   (fifo_empty),
        .fifo_clear   (adc_trig)  // Clear FIFO when ADC is triggered
    );

    // --------------------------------------------------------------------------
    // APB Read
    // --------------------------------------------------------------------------
    // When read enabled, return status register or FIFO data based on address
    always @(posedge PCLK or negedge PRESETn) begin
        if (!PRESETn)
            PRDATA <= 32'b0;
        else if (read_enable) begin
            case (PADDR)
                STATUS_REG_ADDR:     PRDATA <= status_reg;
                MEASUREMENT_HI_ADDR: PRDATA <= fifo_data_out[55:24];
                MEASUREMENT_LO_ADDR: PRDATA <= {8'b0, fifo_data_out[23:0]};
                default:             PRDATA <= 32'b0;
            endcase
        end
        else
            PRDATA <= 32'b0;
    end

    // --------------------------------------------------------------------------
    // The logic for generating the FIFO d_en pulse: When the APB read address is 12'h003 and the FIFO is not empty, 
    // a one cycle high pulse is generated
    // --------------------------------------------------------------------------
    always @(posedge PCLK or negedge PRESETn) begin
        if (!PRESETn)
            fifo_rd_en <= 1'b0;
        else begin
            if (read_enable && (PADDR == MEASUREMENT_LO_ADDR) && !fifo_empty)
                fifo_rd_en <= 1'b1;
            else
                fifo_rd_en <= 1'b0;
        end
    end

    // --------------------------------------------------------------------------
    // Generate a delay signal (delayed by one clock cycle for status updates)
    // --------------------------------------------------------------------------
    always @(posedge PCLK or negedge PRESETn) begin
        if (!PRESETn)
            fifo_rd_en_d <= 1'b0;
        else
            fifo_rd_en_d <= fifo_rd_en;
    end

    // --------------------------------------------------------------------------
    // Status register update: reflects FIFO status and ADC data validity
    // Use the delay signal Fiforud_en-d to determine if a departure has just occurred
    // --------------------------------------------------------------------------
    always @(posedge PCLK or negedge PRESETn) begin
        if (!PRESETn) begin
            status_reg <= 32'b0;
        end else begin
            if (fifo_rd_en_d)
                status_reg[1:0] <= fifo_empty ? 2'b00 : 2'b01;
            else
                status_reg[1:0] <= fifo_empty ? 2'b00 : (fifo_full ? 2'b10 : 2'b01);
            status_reg[3:2] <= adc_data_valid ? 2'b01 : 2'b00;
            status_reg[31:4] <= 28'b0;
        end
    end

    // --------------------------------------------------------------------------
    // APB write operation: Write to PLL, AMUX, and ADC trigger registers
    // --------------------------------------------------------------------------
    // PLL control writing
    always @(posedge PCLK or negedge PRESETn) begin
        if (!PRESETn)
            pll_reg <= {DATA_WIDTH{1'b0}};
        else if (write_enable && (PADDR == PLL_CONTROL_ADDR))
            pll_reg <= PWDATA;
    end

    // AMUX Control Write
    always @(posedge PCLK or negedge PRESETn) begin
        if (!PRESETn)
            amux_reg <= {DATA_WIDTH{1'b0}};
        else if (write_enable && (PADDR == AMUX_ADDR))
            amux_reg <= PWDATA;
    end

    // ADC triggered write: triggered when APB write address is 12'h102,
    // Simultaneously update the trigger register and generate a FIFO reset pulse (adc_rig)
    always @(posedge PCLK or negedge PRESETn) begin
        if (!PRESETn) begin
            trig_reg <= {DATA_WIDTH{1'b0}};
            adc_trig <= 1'b0;
        end else begin
            if (write_enable && (PADDR == ADC_TRIGGER_ADDR)) begin
                trig_reg <= PWDATA;
                adc_trig <= PWDATA[0]; // Use the lowest bit as the trigger signal
            end else begin
                adc_trig <= 1'b0;
            end
        end
    end

    // --------------------------------------------------------------------------
    // APB response logic: Always ready for transmission, no errors occur
    // --------------------------------------------------------------------------
    always @(posedge PCLK) begin
        PREADY <= 1'b1;
    end
    assign PSLVERR = 1'b0;

    // --------------------------------------------------------------------------
    // Debug Output
    // --------------------------------------------------------------------------
    always @(posedge PCLK) begin
        // Debug output can be used to validate write operations 
        // if (write_enable && (PADDR == PLL_CONTROL_ADDR))
        //     $display("PLL_CONTROL: %h", pll_reg);
        // if (write_enable && (PADDR == AMUX_ADDR))
        //     $display("AMUX: %h", amux_reg);
        // if (write_enable && (PADDR == ADC_TRIGGER_ADDR))
        //     $display("ADC_TRIGGER: %h", trig_reg);
    end

    // --------------------------------------------------------------------------
    // INSERT ADC module here.
    // --------------------------------------------------------------------------
    // Dummy ADC 和 AMUX instance
    wire analog_passthrough;
    dummy_adc adc_inst (
        .STATUS_REG_ADDR(status_reg),
        .MEASUREMENT    (fifo_data_out[55:24]), // Retrieve high 32-bit ADC data from FIFO
        .PLL_CONTROL    (pll_reg),
        .ADC_TRIGGER    (trig_reg), 
        .ANALOG_IN      (analog_passthrough)
    );

    dummy_amux amux_inst (
        .INPUT_SEL          (amux_reg[1:0]), 
        .ANALOG_PASSTHROUGH (analog_passthrough)
    );

endmodule
